module lib

pub fn ref[T](v T) &T {
	return &v
}
